LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY encoder2_4 IS
	PORT(w: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		I: OUT STD_LOGIC_VECTOR(3 DOWNTO O));
END decoder2_4;
ARCHITECTURE Behavior OF decoder2_4 IS
BEGIN
	PROCESS(w)
	BEGIN
	CASE w IS
	WHEN "00"=>I<="0000";
	WHEN "01"=>I<="0010";
	WHEN "10"=>I<="0001";
	WHEN "11"=>I<="0101";
	WHEN OTHER =>I<= "XXXX";
	END CASE;
	END PROCESS;
END Behavior;
